module test;

reg clk;
reg [3:0] KEY;
wire [9:0] LEDR;
wire [6:0] HEX5, HEX4, HEX3, HEX2, HEX1, HEX0;

lab1 dut(clk, KEY, LEDR, HEX5, HEX4, HEX3, HEX2, HEX1, HEX0);


  initial begin 
    clk = 1;#10;
    forever begin
      clk = 0; #10;
      clk = 1; #10;
    end
  end

  initial begin 
    KEY = 4'b1111;
    KEY[3] = 1;#10;
    KEY[3] = 0;#10;
    KEY[3] = 1;

    KEY[0] = 1;#50;
    KEY[0] = 0;#10;
    KEY[0] = 1;#100;

    KEY[0] = 0;#10;
    KEY[0] = 1;#100;

    KEY[0] = 0;#10;
    KEY[0] = 1;#100;

    KEY[0] = 0;#10;
    KEY[0] = 1;#100;

    KEY[0] = 0;#10;
    KEY[0] = 1;#100;

    KEY[0] = 0;#10;
    KEY[0] = 1;#100;

    KEY[3] = 1;#10;
    KEY[3] = 0;#10;
    KEY[3] = 1;
    #30;
    KEY[0] = 0;#10;
    KEY[0] = 1;#130;

    KEY[0] = 0;#10;
    KEY[0] = 1;#148;

    KEY[0] = 0;#10;
    KEY[0] = 1;#97;

    KEY[0] = 0;#10;
    KEY[0] = 1;#105;

    KEY[0] = 0;#10;
    KEY[0] = 1;#156;

    KEY[0] = 0;#10;
    KEY[0] = 1;#180;

    KEY[0] = 0;#10;
    KEY[0] = 1;#100;

    KEY[0] = 0;#10;
    KEY[0] = 1;#100;

    
    KEY[0] = 0;#10;
    KEY[0] = 1;#100;
  end

  initial begin
  #150;
    $stop;
  end
endmodule
