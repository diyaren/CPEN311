// Implements a simple Nios II system for the DE-series board.// Inputs:  SW7−0 are parallel port inputs to the Nios II system
//          CLOCK_50 is the system clock
//          KEY[0] is the active-low system reset  // Outputs: LEDR7−0 are parallel port outputs from the Nios II system
module lights (CLOCK_50, SW, KEY, LEDR, HEX1, HEX0, HEX4);input CLOCK_50; 
input [7:0] SW; 
input [0:0] KEY; 
output [7:0] LEDR;output [6:0] HEX1, HEX0, HEX4;wire[7:0] ledConnect;
wire[7:0] prime;// Instantiate the Nios II system module generated by the Qsys tool: 

nios_system NiosII (   .clk_clk(CLOCK_50),    .leddriver1_export(ledConnect),   .prime_export(prime),   .switches_export(SW),    .reset_reset_n(KEY),
   .leds_export(LEDR));

card7seg lightsUp (ledConnect[3:0],HEX0);
card7seg lightsDown(ledConnect[7:4],HEX1);   primeNum primenum(prime[0], HEX4);
	
	endmodule
