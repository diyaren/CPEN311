	component nios_system is
		port (
			clk_clk           : in  std_logic                    := 'X';             -- clk
			leddriver1_export : out std_logic_vector(7 downto 0);                    -- export
			leds_export       : out std_logic_vector(7 downto 0);                    -- export
			reset_reset_n     : in  std_logic                    := 'X';             -- reset_n
			switches_export   : in  std_logic_vector(7 downto 0) := (others => 'X'); -- export
			prime_export      : out std_logic_vector(7 downto 0)                     -- export
		);
	end component nios_system;

	u0 : component nios_system
		port map (
			clk_clk           => CONNECTED_TO_clk_clk,           --        clk.clk
			leddriver1_export => CONNECTED_TO_leddriver1_export, -- leddriver1.export
			leds_export       => CONNECTED_TO_leds_export,       --       leds.export
			reset_reset_n     => CONNECTED_TO_reset_reset_n,     --      reset.reset_n
			switches_export   => CONNECTED_TO_switches_export,   --   switches.export
			prime_export      => CONNECTED_TO_prime_export       --      prime.export
		);

